----------------------------------------------------------------------------------
-- Company:  NIIT University
-- Engineer: Sudhanshu Gupta
-- 
-- Create Date:    16:48:43 10/31/2017
-- Module Name:    gpio_block - Behavioral 
-- Project Name:   processor
-- Target Devices: Numato MIMAS V2
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity gpio_block is
    Port ( DATA_IN   : in    STD_LOGIC_VECTOR (7 downto 0);
           DATA_LOAD : in    STD_LOGIC;
           DIR_LOAD  : in    STD_LOGIC;
           CLOCK     : in    STD_LOGIC;
           DATA_OUT  : out   STD_LOGIC_VECTOR (7 downto 0);
           GPIO      : inout STD_LOGIC_VECTOR (7 downto 0));
end gpio_block;

architecture Behavioral of gpio_block is

   -- import 8-bit register
   component reg8
    Port ( DATA     : in  STD_LOGIC_VECTOR (7 downto 0);
           LOAD_EN  : in  STD_LOGIC;
           RESET    : in  STD_LOGIC;
           CLOCK    : in  STD_LOGIC;
           Q        : out STD_LOGIC_VECTOR (7 downto 0));
   end component;
   
   -- import tristate buffer
   component tristate_buffer
    Port ( A : in  STD_LOGIC;
           G : in  STD_LOGIC;
           Y : out STD_LOGIC);
   end component;
   
   -- direction register signals
   signal DIR_REG_OUT : STD_LOGIC_VECTOR (7 DOWNTO 0);
   
   -- data register signals
   signal DATA_REG_IN : STD_LOGIC_VECTOR (7 DOWNTO 0);
   signal DATA_REG_OUT : STD_LOGIC_VECTOR (7 DOWNTO 0);
   signal DATA_REG_LOAD : STD_LOGIC_VECTOR (7 DOWNTO 0);

begin

   -------------------------
   -- 8 MUXs for DATA_REG_IN
   -------------------------
   with (DIR_REG_OUT(0)) select
      DATA_REG_IN(0) <= GPIO(0)    when '0',
                        DATA_IN(0) when '1',
                        '0'        when others;
   with (DIR_REG_OUT(1)) select
      DATA_REG_IN(1) <= GPIO(1)    when '0',
                        DATA_IN(1) when '1',
                        '0'        when others;
   with (DIR_REG_OUT(2)) select
      DATA_REG_IN(2) <= GPIO(2)    when '0',
                        DATA_IN(2) when '1',
                        '0'        when others;
   with (DIR_REG_OUT(3)) select
      DATA_REG_IN(3) <= GPIO(3)    when '0',
                        DATA_IN(3) when '1',
                        '0'        when others;
   with (DIR_REG_OUT(4)) select
      DATA_REG_IN(4) <= GPIO(4)    when '0',
                        DATA_IN(4) when '1',
                        '0'        when others;
   with (DIR_REG_OUT(5)) select
      DATA_REG_IN(5) <= GPIO(5)    when '0',
                        DATA_IN(5) when '1',
                        '0'        when others;
   with (DIR_REG_OUT(6)) select
      DATA_REG_IN(6) <= GPIO(6)    when '0',
                        DATA_IN(6) when '1',
                        '0'        when others;
   with (DIR_REG_OUT(7)) select
      DATA_REG_IN(7) <= GPIO(7)    when '0',
                        DATA_IN(7) when '1',
                        '0'        when others;
   
   ---------------------------
   -- 8 MUXs for DATA_REG_LOAD
   ---------------------------
   with (DIR_REG_OUT(0)) select
      DATA_REG_LOAD(0) <= '1'       when '0',
                          DATA_LOAD when '1',
                          '0'       when others;
   with (DIR_REG_OUT(1)) select
      DATA_REG_LOAD(1) <= '1'       when '0',
                          DATA_LOAD when '1',
                          '0'       when others;
   with (DIR_REG_OUT(2)) select
      DATA_REG_LOAD(2) <= '1'       when '0',
                          DATA_LOAD when '1',
                          '0'       when others;
   with (DIR_REG_OUT(3)) select
      DATA_REG_LOAD(3) <= '1'       when '0',
                          DATA_LOAD when '1',
                          '0'       when others;
   with (DIR_REG_OUT(4)) select
      DATA_REG_LOAD(4) <= '1'       when '0',
                          DATA_LOAD when '1',
                          '0'       when others;
   with (DIR_REG_OUT(5)) select
      DATA_REG_LOAD(5) <= '1'       when '0',
                          DATA_LOAD when '1',
                          '0'       when others;
   with (DIR_REG_OUT(6)) select
      DATA_REG_LOAD(6) <= '1'       when '0',
                          DATA_LOAD when '1',
                          '0'       when others;
   with (DIR_REG_OUT(7)) select
      DATA_REG_LOAD(7) <= '1'       when '0',
                          DATA_LOAD when '1',
                          '0'       when others;
   
   DATA_OUT <= DATA_REG_OUT;

   -- 8-bit data register, with separate LOAD for each bit
   data_reg_inst: process(CLOCK)
   begin
      if (rising_edge(CLOCK)) then
         if (DATA_REG_LOAD(0) = '1') then
            DATA_REG_OUT(0) <= DATA_REG_IN(0);
         end if;
         if (DATA_REG_LOAD(1) = '1') then
            DATA_REG_OUT(1) <= DATA_REG_IN(1);
         end if;
         if (DATA_REG_LOAD(2) = '1') then
            DATA_REG_OUT(2) <= DATA_REG_IN(2);
         end if;
         if (DATA_REG_LOAD(3) = '1') then
            DATA_REG_OUT(3) <= DATA_REG_IN(3);
         end if;
         if (DATA_REG_LOAD(4) = '1') then
            DATA_REG_OUT(4) <= DATA_REG_IN(4);
         end if;
         if (DATA_REG_LOAD(5) = '1') then
            DATA_REG_OUT(5) <= DATA_REG_IN(5);
         end if;
         if (DATA_REG_LOAD(6) = '1') then
            DATA_REG_OUT(6) <= DATA_REG_IN(6);
         end if;
         if (DATA_REG_LOAD(7) = '1') then
            DATA_REG_OUT(7) <= DATA_REG_IN(7);
         end if;
      end if;
   end process data_reg_inst;
   
   -- 8-bit direction register
   dir_reg_inst: reg8
      PORT MAP (
         DATA => DATA_IN,
         LOAD_EN => DIR_LOAD,
         RESET => '0',
         CLOCK => CLOCK,
         Q => DIR_REG_OUT
      );
   
   -----------------------------------------------
   -- 8 tristate buffers to control output to GPIO
   -----------------------------------------------
   tsb0: tristate_buffer
      PORT MAP (
         A => DATA_REG_OUT(0),
         G => DIR_REG_OUT(0),
         Y => GPIO(0)
      );
   tsb1: tristate_buffer
      PORT MAP (
         A => DATA_REG_OUT(1),
         G => DIR_REG_OUT(1),
         Y => GPIO(1)
      );
   tsb2: tristate_buffer
      PORT MAP (
         A => DATA_REG_OUT(2),
         G => DIR_REG_OUT(2),
         Y => GPIO(2)
      );
   tsb3: tristate_buffer
      PORT MAP (
         A => DATA_REG_OUT(3),
         G => DIR_REG_OUT(3),
         Y => GPIO(3)
      );
   tsb4: tristate_buffer
      PORT MAP (
         A => DATA_REG_OUT(4),
         G => DIR_REG_OUT(4),
         Y => GPIO(4)
      );
   tsb5: tristate_buffer
      PORT MAP (
         A => DATA_REG_OUT(5),
         G => DIR_REG_OUT(5),
         Y => GPIO(5)
      );
   tsb6: tristate_buffer
      PORT MAP (
         A => DATA_REG_OUT(6),
         G => DIR_REG_OUT(6),
         Y => GPIO(6)
      );
   tsb7: tristate_buffer
      PORT MAP (
         A => DATA_REG_OUT(7),
         G => DIR_REG_OUT(7),
         Y => GPIO(7)
      );

end Behavioral;
